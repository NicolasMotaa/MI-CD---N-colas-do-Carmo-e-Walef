module subtrator4x4 (S, Bo, A, B, Bin);

    input [3:0] A, B; 
    input Bin; 
    output [3:0] S;
    output Bo;

    wire c1, c2, c3;

    // Instanciando o subtrator de 1 bit para cada bit
    subtratorbase s0 (.A(A[0]), .B(B[0]), .Bin(Bin),  .S(S[0]), .Bo(c1));
    subtratorbase s1 (.A(A[1]), .B(B[1]), .Bin(c1),   .S(S[1]), .Bo(c2));
    subtratorbase s2 (.A(A[2]), .B(B[2]), .Bin(c2),   .S(S[2]), .Bo(c3));
    subtratorbase s3 (.A(A[3]), .B(B[3]), .Bin(c3),   .S(S[3]), .Bo(Bo));

endmodule